module multi_fix #(parameter WORDLENGTH = 8, FRACTION = 4)(
  output signed

)
