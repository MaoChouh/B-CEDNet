/*
    Copyright
    All right reserved.
    Author  : Zichuan Liu, Yixing Li and Wenye Liu.
    Description: This is the global parameters file that configures the architecture of the design.
*/


`define MODE_SIM