/*
Copyright
All right reserved.
Author  : Zichuan Liu, Yixing Li and Wenye Liu.
Description: This is the header file for configure the testbench_PE_FP.
*/

`define PARAM_INPUTPATH "../../test/testbench_PE_FP/input/"
`define PARAM_OUTPUTPATH "../../test/testbench_PE_FP/output/"
`define PARAM_TESTBENCH testbench_PE_FP
`define PARAM_D 1
`define PARAM_FH 3
`define PARAM_FW 3
`define PARAM_POOL_H 1
`define PARAM_POOL_W 1
`define PARAM_STRIDE_H 1
`define PARAM_STRIDE_W 1
`define PARAM_DATA_IN_FP_WIDTH 17
`define PARAM_DATA_IN_FP_FRAC_WIDTH 8
`define PARAM_WEIGHT_WIDTH 17
`define PARAM_WEIGHT_FRAC_WIDTH 8
`define PARAM_IN_WINDOW_H 3
`define PARAM_IN_WINDOW_W 3
`define PARAM_REF_WIDTH 22
`define PARAM_IN_WIDTH 153
`define PARAM_OUT_WIDTH 1
