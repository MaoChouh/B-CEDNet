/*
Copyright
All right reserved.
Author  : Zichuan Liu, Yixing Li and Wenye Liu.
Description: This is the header file for configure the TOP.
*/

`define PARAM_TOP_INPUTPATH "../../test/TOP/input/"
`define PARAM_TOP_OUTPUTPATH "../../test/TOP/output/"
`define PARAM_TOP_BLOCK_NAME TOP
`define PARAM_TOP_MEAN_ROM_NAME "TOP_MEAN_ROM"
`define PARAM_TOP_MEAN_WIDTH 17
`define PARAM_TOP_MEAN_FRAC_WIDTH 8
`define PARAM_TOP_MEAN_ROM_DEPTH 4096
`define PARAM_TOP_MEAN_ROM_INST_TYPE "FULL_SOFT"
