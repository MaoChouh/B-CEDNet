/*
Copyright
All right reserved.
Author  : Zichuan Liu, Yixing Li and Wenye Liu.
Description: This is the header file for configure the ROM_SOFT_F_tb.
*/

`define PARAM_INPUTPATH "../../test/ROM_SOFT_F_tb/input/"
`define PARAM_OUTPUTPATH "../../test/ROM_SOFT_F_tb/output/"
`define PARAM_TESTBENCH ROM_SOFT_F_tb
`define PARAM_DATA_WIDTH 4608
`define PARAM_DATA_DEPTH 64
`define PARAM_DATA_DIV 12
`define PARAM_CLK_PERIOD 130
`define PARAM_CLK_R_PERIOD 10
`define PARAM_TRUE_DATA_WITH 384
`define PARAM_TRUE_DATA_DEPTH 768
`define PARAM_ROM_NAME "ROM_CORE_TEST"
