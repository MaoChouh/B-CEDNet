/*
Copyright
All right reserved.
Author  : Zichuan Liu, Yixing Li and Wenye Liu.
Description: This is the header file for configure the W_ROM_tb.
*/

`define PARAM_INPUTPATH "../../test/W_ROM_tb/input/"
`define PARAM_OUTPUTPATH "../../test/W_ROM_tb/output/"
`define PARAM_TESTBENCH W_ROM_tb
`define PARAM_DATA_WIDTH 1152
`define PARAM_DATA_DEPTH 128
`define PARAM_INST_TYPE "FULL_SOFT"
`define PARAM_PRELOADFILE ""
`define PARAM_ADDR_WIDTH 7
`define PARAM_CLK_PERIOD 10
`define PARAM_MEM_NAME "W_ROM_SOFT_T"
