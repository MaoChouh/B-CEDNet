/*
Copyright
All right reserved.
Author  : Zichuan Liu, Yixing Li and Wenye Liu.
Description: This is the header file for configure the testbench_PE_DC.
*/

`define PARAM_INPUTPATH "../../test/testbench_PE_DC/input/"
`define PARAM_OUTPUTPATH "../../test/testbench_PE_DC/output/"
`define PARAM_TESTBENCH testbench_PE_DC
`define PARAM_D 512
`define PARAM_FH 3
`define PARAM_FW 3
`define PARAM_POOL_H 2
`define PARAM_POOL_W 2
`define PARAM_STRIDE_H 1
`define PARAM_STRIDE_W 1
`define PARAM_REF_WIDTH 14
`define PARAM_PINDEX_WIDTH 2
`define PARAM_IN_WIDTH 4608
`define PARAM_OUT_WIDTH 4
