/*
Copyright
All right reserved.
Author  : Zichuan Liu, Yixing Li and Wenye Liu.
Description: This is the header file for configure the BCEDN_TOP_tb.
*/

`define PARAM_INPUTPATH "F:/Vivado_prj/B-CEDNet/test/BCEDN_TOP_tb/input/"
`define PARAM_OUTPUTPATH "F:/Vivado_prj/B-CEDNet/test/BCEDN_TOP_tb/output/"
`define PARAM_TESTBENCH BCEDN_TOP_tb
`define PARAM_DATA_IN_WIDTH 8
`define PARAM_CLK_DIV 13
`define PARAM_DATA_OUT_WIDTH 24
`define PARAM_CLK_P_PERIOD 130
`define PARAM_CLK_R_PERIOD 10
`define PARAM_PROCESSING_CYC 786432
