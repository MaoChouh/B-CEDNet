`define LOAD_MEM initial begin \
if (INST_TYPE != "FULL_SOFT") begin\
end\
end
