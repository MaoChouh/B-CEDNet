/*
Copyright
All right reserved.
Author  : Zichuan Liu, Yixing Li and Wenye Liu.
Description: This is the header file for configure the testbench_PE_EC.
*/

`define PARAM_INPUTPATH "F:/Vivado_prj/B-CEDNet/test/testbench_PE_EC/input/"
`define PARAM_OUTPUTPATH "F:/Vivado_prj/B-CEDNet/test/testbench_PE_EC/output/"
`define PARAM_TESTBENCH testbench_PE_EC
`define PARAM_D 128
`define PARAM_FH 3
`define PARAM_FW 3
`define PARAM_POOL_H 2
`define PARAM_POOL_W 2
`define PARAM_STRIDE_H 1
`define PARAM_STRIDE_W 1
`define PARAM_IN_WINDOW_H 4
`define PARAM_IN_WINDOW_W 4
`define PARAM_REF_WIDTH 12
`define PARAM_IN_WIDTH 2048
`define PARAM_PINDEX_WIDTH 2
`define PARAM_OUT_WIDTH 1
