/*
Copyright
All right reserved.
Author  : Zichuan Liu, Yixing Li and Wenye Liu.
Description: This is the header file for configure the DC_10.
*/

`define PARAM_DC_10_INPUTPATH "../../test/DC_10/input/"
`define PARAM_DC_10_OUTPUTPATH "../../test/DC_10/output/"
`define PARAM_DC_10_BLOCK_NAME DC_10
`define PARAM_DC_10_M 1
`define PARAM_DC_10_P 1
`define PARAM_DC_10_H 128
`define PARAM_DC_10_W 32
`define PARAM_DC_10_D 512
`define PARAM_DC_10_FH 1
`define PARAM_DC_10_FW 1
`define PARAM_DC_10_FD 27
`define PARAM_DC_10_PAD 1
`define PARAM_DC_10_STRIDE_H 1
`define PARAM_DC_10_STRIDE_W 1
`define PARAM_DC_10_POOL_H 1
`define PARAM_DC_10_POOL_W 1
`define PARAM_DC_10_N_PE 1
`define PARAM_DC_10_NORMREF_SCALE_WIDTH 12
`define PARAM_DC_10_NORMREF_SCALE_FRAC_WIDTH 11
`define PARAM_DC_10_REF_WIDTH_FROM_NET 8
`define PARAM_DC_10_NORMREF_WIDTH 12
`define PARAM_DC_10_DATA_OUT_WIDTH 24
`define PARAM_DC_10_ROM_INST_TYPE "FULL_SOFT"
`define PARAM_DC_10_W_MEM_NAME "DC_10_W_ROM"
`define PARAM_DC_10_REF_MEM_NAME "DC_10_REF_ROM"
`define PARAM_DC_10_REF_SCALE_MEM_NAME "DC_10_REF_SCALE_ROM"
`define PARAM_DC_10_ROM_INDEX {0}
